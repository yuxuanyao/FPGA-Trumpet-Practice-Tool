
module AudioV2 (
	// Inputs
	CLOCK_50,
	KEY,

	AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	FPGA_I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,

	FPGA_I2C_SCLK,
	SW
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input				CLOCK_50;
input		[3:0]	KEY;
input		[3:0]	SW;

input				AUD_ADCDAT;

// Bidirectionals
inout				AUD_BCLK;
inout				AUD_ADCLRCK;
inout				AUD_DACLRCK;

inout				FPGA_I2C_SDAT;

// Outputs
output				AUD_XCK;
output				AUD_DACDAT;

output				FPGA_I2C_SCLK;

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
// Internal Wires
wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
wire				read_audio_in;

wire				audio_out_allowed;
wire		[31:0]	left_channel_audio_out;
wire		[31:0]	right_channel_audio_out;
wire				write_audio_out;

wire resetcounter;
assign resetcounter = KEY[1];

// Internal Registers


reg [14:0] delay_cnt;
wire [14:0] delay;
reg [15:0] m;
reg [15:0] rate = 16'd 5000;
reg [15:0] counter ;
reg [15:0] a;
reg snd;

reg [8:0] cnt ;
wire [15:0] count = 16'd2000;

wire [5:0] audio_from_ram;
wire [13:0] address_count;

reg [13:0] address_count_reg;
reg [10:0] clk_count;


ram_1 memory1(
.address(address_count),
.clock(CLOCK_50),
.data(),
.wren(1'b0),
.q(audio_from_ram));


// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/


/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/
always @(posedge CLOCK_50)begin
	if(clk_count == 11'd1200)  begin
		if(address_count_reg == 14'd16383) begin
			address_count_reg <= 14'b0;
		end 
	else address_count_reg <= address_count_reg + 1;
	clk_count <= 0;
	
end 
else
	clk_count <= clk_count + 1;
end
assign address_count = address_count_reg;
	
	/*
	if (!resetcounter) begin
		m <= 16'd0;
		counter <= 16'd0;
		end
	else if (counter == rate) begin
		m <= m + 1;
		counter <= 16'd0;
		end
	else
		counter <= counter + 1;
  */
 
/* always @(m)
	 begin
	 if ( m < count)
		a <= m;
		else
		m <= 16'd0;
	end */
 
/*always @(m)
	if(delay_cnt == delay) begin
		delay_cnt <= 0;
		snd <= !snd;
	end else delay_cnt <= delay_cnt + 1;*/

/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/

assign delay = {15'd100};

//wire [31:0] sound = (SW == 0) ? 0 : snd ? 32'd10000000 : -32'd10000000;


assign read_audio_in			= audio_in_available & audio_out_allowed;

assign left_channel_audio_out	= {audio_from_ram, 26'b0};
assign right_channel_audio_out	= 32'b0;

assign write_audio_out			= audio_in_available & audio_out_allowed;

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

Audio_Controller Audio_Controller (
	// Inputs
	.CLOCK_50						(CLOCK_50),
	.reset						(~KEY[0]),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out ),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),


	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)

);

avconf #(.USE_MIC_INPUT(1)) avc (
	.FPGA_I2C_SCLK					(FPGA_I2C_SCLK),
	.FPGA_I2C_SDAT					(FPGA_I2C_SDAT),
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0])
);

endmodule

